	package enum_pkg;
		typedef enum logic [1:0] {
			NO_PARITY 	= 2'b00,
			ODD_PARITY 	= 2'b01,
			EVEN_PARITY = 2'b10
		} parity_t;
		
	endpackage : enum_pkg
